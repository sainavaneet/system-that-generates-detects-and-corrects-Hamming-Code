`timescale 1ns / 1ps

module hamming_tb();

reg [6:0] part_7790_0, part_7790_1, part_7790_2, part_7790_3, part_7790_4, part_7790_5, part_7790_6, 
          part_7790_7, part_7790_8, part_7790_9, part_7790_10, part_7790_11, part_7790_12, 
          part_7790_13, part_7790_14, part_7790_15;

wire [10:0] out_77990_0, out_77990_1, out_77990_2, out_77990_3, out_77990_4, out_77990_5, out_77990_6, out_77990_7, out_77990_8, out_77990_9, out_77990_10, out_77990_11, 
            out_77990_12, out_77990_13, out_77990_14, out_77990_15;

hamming hu(.part_7790_0(part_7790_0), .part_7790_1(part_7790_1), 
            .part_7790_2(part_7790_2), .part_7790_3(part_7790_3), 
            .part_7790_4(part_7790_4), .part_7790_5(part_7790_5), 
            .part_7790_6(part_7790_6), .part_7790_7(part_7790_7), 
            .part_7790_8(part_7790_8), .part_7790_9(part_7790_9), 
            .part_7790_10(part_7790_10), .part_7790_11(part_7790_11), 
            .part_7790_12(part_7790_12), .part_7790_13(part_7790_13), 
            .part_7790_14(part_7790_14), .part_7790_15(part_7790_15),
            .out_77990_0(out_77990_0), .out_77990_1(out_77990_1), .out_77990_2(out_77990_2), .out_77990_3(out_77990_3), .out_77990_4(out_77990_4), .out_77990_5(out_77990_5), 
            .out_77990_6(out_77990_6), .out_77990_7(out_77990_7), .out_77990_8(out_77990_8), .out_77990_9(out_77990_9), .out_77990_10(out_77990_10), .out_77990_11(out_77990_11), 
            .out_77990_12(out_77990_12), .out_77990_13(out_77990_13), .out_77990_14(out_77990_14), .out_77990_15(out_77990_15));




initial begin

    part_7790_0 = 7'b1001000;
    #2;
    part_7790_1 = 7'b1100101;
    #2;
    part_7790_2 = 7'b1101100;
    #2;
    part_7790_3 = 7'b1101100;
    #2;
    part_7790_4 = 7'b1101111;
    #2;
    part_7790_5 = 7'b0100000;
    #2;
    part_7790_6 = 7'b1000011;
    #2;
    part_7790_7 = 7'b1001111;
    #2;
    part_7790_8 = 7'b1001101;
    #2;
    part_7790_9 = 7'b1010000;
    #2;
    part_7790_10 = 7'b0110011;
    #2;
    part_7790_11 = 7'b0110001;
    #2;
    part_7790_12 = 7'b0110001;
    #2;
    part_7790_13 = 7'b0101101;
    #2;
    part_7790_14 = 7'b0110010;
    #2;
    part_7790_15 = 7'b0100001;
    #2;


   $display("--------------------------------------------------------------------");


    $display("out_77990_0  = %h", out_77990_0);
    $display("out_77990_1  = %h", out_77990_1);
    $display("out_77990_2  = %h", out_77990_2);
    $display("out_77990_3  = %h", out_77990_3);
    $display("out_77990_4  = %h", out_77990_4);
    $display("out_77990_5  = %h", out_77990_5);
    $display("out_77990_6  = %h", out_77990_6);
    $display("out_77990_7  = %h", out_77990_7);
    $display("out_77990_8  = %h", out_77990_8);
    $display("out_77990_9  = %h", out_77990_9);
    $display("out_77990_10 = %h", out_77990_10);
    $display("out_77990_11 = %h", out_77990_11);
    $display("out_77990_12 = %h", out_77990_12);
    $display("out_77990_13 = %h", out_77990_13);
    $display("out_77990_14 = %h", out_77990_14);
    $display("out_77990_15 = %h", out_77990_15);

end






    
endmodule